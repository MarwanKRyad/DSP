module DSP_tb();

reg [17:0] A,B,D;
reg [47:0] C;
reg clk,CARRYIN;
reg [7:0] OPMODE;
reg [17:0] BCIN;
reg RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE;
reg [47:0]PCIN ;
wire [17:0]BCOUT;
wire [47:0]PCOUT;
wire [47:0]P;
wire [35:0]M;
wire CARRYOUT;
wire CARRYOUTF;
DSP DUT(A,B,C,D,clk,CARRYIN,OPMODE,BCIN,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE,PCIN,BCOUT,PCOUT,P,M,CARRYOUT,CARRYOUTF);

initial begin
	clk=0;
	forever 
	#1 clk=~clk;		
end
initial
begin

A=1;B=1;C=1;D=1;CARRYIN=1;OPMODE=8'b01111101;BCIN=0;RSTA=0;RSTB=0;RSTM=0;RSTP=0;RSTC=0;RSTD=0;RSTCARRYIN=0;RSTOPMODE=0;
CEA=1;CEB=1;CEM=1;CEP=1;CEC=1;CED=1;CECARRYIN=1;CEOPMODE=1;PCIN=0;
//p=[(B-D)*A+opmode[5]+c]=2
#8
A=1;B=1;C=1;D=1;CARRYIN=1;OPMODE=8'b00111101;BCIN=0;RSTA=0;RSTB=0;RSTM=0;RSTP=0;RSTC=0;RSTD=0;RSTCARRYIN=0;RSTOPMODE=0;
CEA=1;CEB=1;CEM=1;CEP=1;CEC=1;CED=1;CECARRYIN=1;CEOPMODE=1;PCIN=0;
//p=[(B+D)*A+opmode[5]+c]=4


#8

A=1;B=1;C=3;D=1;CARRYIN=1;OPMODE=8'b00011101;BCIN=0;RSTA=0;RSTB=0;RSTM=0;RSTP=0;RSTC=0;RSTD=0;RSTCARRYIN=0;RSTOPMODE=0;
CEA=1;CEB=1;CEM=1;CEP=1;CEC=1;CED=1;CECARRYIN=1;CEOPMODE=1;PCIN=0;
//p=[(B+D)*A+c]=5
#8

A=1;B=1;C=3;D=1;CARRYIN=1;OPMODE=8'b00111100;BCIN=0;RSTA=0;RSTB=0;RSTM=0;RSTP=0;RSTC=0;RSTD=0;RSTCARRYIN=0;RSTOPMODE=0;
CEA=1;CEB=1;CEM=1;CEP=1;CEC=1;CED=1;CECARRYIN=1;CEOPMODE=1;PCIN=0;
//p=c+opmode[5]=4

#8
A=1;B=1;C=3;D=1;CARRYIN=1;OPMODE=8'b00110000;BCIN=0;RSTA=0;RSTB=0;RSTM=0;RSTP=0;RSTC=0;RSTD=0;RSTCARRYIN=0;RSTOPMODE=0;
CEA=1;CEB=1;CEM=1;CEP=1;CEC=1;CED=1;CECARRYIN=1;CEOPMODE=1;PCIN=0;
//p=opmode[5]=1
#8
A=1;B=1;C=3;D=1;CARRYIN=1;OPMODE=8'b00010000;BCIN=0;RSTA=0;RSTB=0;RSTM=0;RSTP=0;RSTC=0;RSTD=0;RSTCARRYIN=0;RSTOPMODE=0;
CEA=1;CEB=1;CEM=1;CEP=1;CEC=1;CED=1;CECARRYIN=1;CEOPMODE=1;PCIN=0;
//p=opmode[5]=0



end
endmodule